module fulladd(input a, input b,input c, output s);

assign s=a^b^c;

endmodule